////////////////////////////////////////////////////////////////////////////////////////////////////
// This program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public License
// as published by the Free Software Foundation; either version 2
// of the License, or (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA
// 02111-1307, USA.
//
// ©2013 - Roman Ovseitsev <romovs@gmail.com>
////////////////////////////////////////////////////////////////////////////////////////////////////

//##################################################################################################
//
// Register configuration for OV7670 camera module.
//
// Initializes RGB565 VGA, with distorted colors... I yet to find the register settings to fix this. 
//
//##################################################################################################

`timescale 1ns / 1ps

module OV7670Init (index_i, data_o);

   input       [5:0] index_i;    // Register index.
   output reg  [16:0] data_o;    // {Register_address, register_value, rw_flag} :
                                 //  Where register_value is the value to write if rw_flag = 1
                                 //  otherwise it's not used when rw_flag = 0 (read).
                                 // {16'hffff, 1'b1} - denotes end of the register set.
                                 // {16'hf0f0, 1'b1} - denotes that a delay is needed at this point.
   always @* begin
      (* parallel_case *) case(index_i)
         //7'd0 : data_o = {16'h0A76, 1'b0}; 
         8'd0 : data_o = {16'h1280, 1'b1};   // COM7     Reset.
         8'd1 : data_o = {16'hf0f0, 1'b1};   // Denotes delay.
         8'd2 : data_o = {16'h1204, 1'b1};   // COM7     Set RGB (06 enables color bar overlay).
         8'd3 : data_o = {16'h1100, 1'b1};   // CLKRC    Use external clock directly.
         8'd4 : data_o = {16'h0C00, 1'b1};   // COM3     Disable DCW & scalling. + RSVD bits.
         8'd5 : data_o = {16'h3E00, 1'b1};   // COM14    Normal PCLK.
         8'd6 : data_o = {16'h8C00, 1'b1};   // RGB444   Disable RGB444
         8'd7 : data_o = {16'h0400, 1'b1};   // COM1     Disable CCIR656. AEC low 2 LSB.
         8'd8 : data_o = {16'h40d0, 1'b1};   // COM15    Set RGB565 full value range
         8'd9 : data_o = {16'h3a04, 1'b1};   // TSLB     Don't set window automatically. + RSVD bits.
         8'd10: data_o = {16'h1418, 1'b1};   // COM9     Maximum AGC value x4. Freeze AGC/AEC. + RSVD bits.
         8'd11: data_o = {16'h4fb3, 1'b1};   // MTX1     Matrix Coefficient 1
         8'd12: data_o = {16'h50b3, 1'b1};   // MTX2     Matrix Coefficient 2
         8'd13: data_o = {16'h5100, 1'b1};   // MTX3     Matrix Coefficient 3
         8'd14: data_o = {16'h523d, 1'b1};   // MTX4     Matrix Coefficient 4
         8'd15: data_o = {16'h53a7, 1'b1};   // MTX5     Matrix Coefficient 5
         8'd16: data_o = {16'h54e4, 1'b1};   // MTX6     Matrix Coefficient 6
         8'd17: data_o = {16'h589e, 1'b1};   // MTXS     Enable auto contrast center. Matrix coefficient sign. + RSVD bits.
         8'd18: data_o = {16'h3dc0, 1'b1};   // COM13    Gamma enable. + RSVD bits.
         8'd19: data_o = {16'h1100, 1'b1};   // CLKRC    Use external clock directly.
         8'd20: data_o = {16'h1714, 1'b1};   // HSTART   HREF start high 8 bits.
         8'd21: data_o = {16'h1802, 1'b1};   // HSTOP    HREF stop high 8 bits.
         8'd22: data_o = {16'h3280, 1'b1};   // HREF     HREF edge offset. HSTART/HSTOP low 3 bits.
         8'd23: data_o = {16'h1903, 1'b1};   // VSTART   VSYNC start high 8 bits.
         8'd24: data_o = {16'h1A7b, 1'b1};   // VSTOP    VSYNC stop high 8 bits.
         8'd25: data_o = {16'h030a, 1'b1};   // VREF     VSYNC edge offset. VSTART/VSTOP low 3 bits.
         8'd26: data_o = {16'h0f41, 1'b1};   // COM6     Disable HREF at optical black. Reset timings. + RSVD bits.
         8'd27: data_o = {16'h1e03, 1'b1};   // MVFP     No mirror/vflip. Black sun disable. + RSVD bits.
         8'd28: data_o = {16'h330b, 1'b1};   // CHLF     Array Current Control - Reserved  
         //8'd29: data_o = {16'h373f, 1'b1};   // ADC 
         //8'd30: data_o = {16'h3871, 1'b1};   // ACOM     ADC and Analog Common Mode Control - Reserved
         //8'd31: data_o = {16'h392a, 1'b1};   // OFON     ADC Offset Control - Reserved               
         8'd29: data_o = {16'h3c78, 1'b1};   // COM12    No HREF when VSYNC is low. + RSVD bits.
         8'd30: data_o = {16'h6900, 1'b1};   // GFIX     Fix Gain Control? No.    
         8'd31: data_o = {16'h6b1a, 1'b1};   // DBLV     Bypass PLL. Enable internal regulator. + RSVD bits.
         8'd32: data_o = {16'h7400, 1'b1};   // REG74    Digital gain controlled by VREF[7:6]. + RSVD bits.
         8'd33: data_o = {16'hb084, 1'b1};   // RSVD     ?          
         8'd34: data_o = {16'hb10c, 1'b1};   // ABLC1    Enable ABLC function. + RSVD bits.
         8'd35: data_o = {16'hb20e, 1'b1};   // RSVD     ?
         8'd36: data_o = {16'hb380, 1'b1};   // THL_ST   ABLC Target.
         /*8'd37: data_o = {16'h7a20, 1'b1};   // SLOP     Gamma Curve Highest Segment Slope 
         8'd38: data_o = {16'h7b10, 1'b1};   // GAM1
         8'd39: data_o = {16'h7c1e, 1'b1};   // GAM2
         8'd40: data_o = {16'h7d35, 1'b1};   // GAM3
         8'd41: data_o = {16'h7e5a, 1'b1};   // GAM4
         8'd42: data_o = {16'h7f69, 1'b1};   // GAM5
         8'd43: data_o = {16'h8076, 1'b1};   // GAM6
         8'd44: data_o = {16'h8180, 1'b1};   // GAM7
         8'd45: data_o = {16'h8288, 1'b1};   // GAM8
         8'd46: data_o = {16'h838f, 1'b1};   // GAM9
         8'd47: data_o = {16'h8496, 1'b1};   // GAM10
         8'd48: data_o = {16'h85a3, 1'b1};   // GAM11
         8'd49: data_o = {16'h86af, 1'b1};   // GAM12
         8'd50: data_o = {16'h87c4, 1'b1};   // GAM13
         8'd51: data_o = {16'h88d7, 1'b1};   // GAM14
         8'd52: data_o = {16'h89e8, 1'b1};   // GAM15*/
         default: data_o = {16'hffff, 1'b1};
      endcase
   end

endmodule
